`include "deco.v"
module top();
  sevenSegmentDecoder_tb UUT();
endmodule
